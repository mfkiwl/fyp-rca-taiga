package rca_config
    localparam NUM_RCAS = 4;
    localparam NUM_READ_PORTS = 5;
    localparam NUM_WRITE_PORTS = 5;


    //RCA Instructions will be of U-type with immediate specifying which accelerator to use (for now) TODO: change to R-type to allow RCA configuration

endpackage