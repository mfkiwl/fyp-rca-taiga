package rca_config
    localparam NUM_RCAS = 4;
    localparam NUM_READ_PORTS = 5;
    localparam NUM_WRITE_PORTS = 5;


    //RCA Instructions will have bits 6:0 as opcode, rest of the bits as accelerator selector 31:7

endpackage